.title KiCad schematic
JB-IN1 Net-_CB1-Pad1_ GND Conn_Coaxial
LB1 Net-_CB1-Pad1_ GND L
CB1 Net-_CB1-Pad1_ GND C
CB2 Net-_CB2-Pad1_ Net-_CB2-Pad2_ C
LB2 Net-_CB1-Pad1_ Net-_CB2-Pad2_ L
JB-OUT1 Net-_CB6-Pad1_ GND Conn_Coaxial
LB3 Net-_CB2-Pad1_ GND L
LB5 Net-_CB4-Pad1_ GND L
CB3 Net-_CB2-Pad1_ GND C
CB5 Net-_CB4-Pad1_ GND C
LB4 Net-_CB2-Pad1_ Net-_CB4-Pad2_ L
CB4 Net-_CB4-Pad1_ Net-_CB4-Pad2_ C
LB6 Net-_CB4-Pad1_ Net-_CB6-Pad2_ L
CB6 Net-_CB6-Pad1_ Net-_CB6-Pad2_ C
JC-IN1 Net-_CC1-Pad1_ GND Conn_Coaxial
CC1 Net-_CC1-Pad1_ GND C
LC1 Net-_CC1-Pad1_ Net-_CC2-Pad1_ L
JC-OUT1 Net-_CC4-Pad1_ GND Conn_Coaxial
CC2 Net-_CC2-Pad1_ GND C
CC3 Net-_CC3-Pad1_ GND C
LC2 Net-_CC2-Pad1_ Net-_CC3-Pad1_ L
LC3 Net-_CC3-Pad1_ Net-_CC4-Pad1_ L
CC4 Net-_CC4-Pad1_ GND C
LB7 Net-_CB6-Pad1_ GND L
CB7 Net-_CB6-Pad1_ GND C
.end
