.MODEL ONSEMI_MMBT5179 NPN (Is=69.28E-18  Xti=3  Eg=1.11  Vaf=100  Bf=282.1  Ne=1.177  Ise=69.28E-18  Ikf=22.03m  Xtb=1.5  Br=1.176 Nc=2    Isc=0    Ikr=0    Rc=4    Cjc=1.042p    Mjc=.2468    Vjc=.75    Fc=.5    Cje=1.52p    Mje=.3223    Vje=.75    Tr=1.588n Tf=135.6p  Itf=.27  Vtf=10  Xtf=30  Rb=10)

.MODEL ONSEMI_2N3904 NPN (IS=1.26532e-10 BF=206.302 NF=1.5 VAF=1000 IKF=0.0272221 ISE=2.30771e-09 NE=3.31052 BR=20.6302 NR=2.89609 VAR=9.39809 IKR=0.272221 ISC=2.30771e-09 NC=1.9876 RB=5.8376 IRB=50.3624 RBM=0.634251 RE=0.0001 RC=2.65711 XTB=0.1 XTI=1 EG=1.05 CJE=4.64214e-12 VJE=0.4 MJE=0.256227 TF=4.19578e-10 XTF=0.906167 VTF=8.75418 ITF=0.0105823 CJC=3.76961e-12 VJC=0.4 MJC=0.238109 XCJC=0.8 FC=0.512134 CJS=0 VJS=0.75 MJS=0.5 TR=6.82023e-08 PTF=0 KF=0 AF=1)

.MODEL ONSEMI_2N2222a NPN (IS=3.88184e-14 BF=929.846 NF=1.10496 VAF=16.5003 IKF=0.019539 ISE=1.0168e-11 NE=1.94752 BR=48.4545 NR=1.07004 VAR=40.538 IKR=0.19539 ISC=1.0168e-11 NC=4 RB=0.1 IRB=0.1 RBM=0.1 RE=0.0001 RC=0.426673 XTB=0.1 XTI=1 EG=1.05 CJE=2.23677e-11 VJE=0.582701 MJE=0.63466 TF=4.06711e-10 XTF=3.92912 VTF=17712.6 ITF=0.4334 CJC=2.23943e-11 VJC=0.576146 MJC=0.632796 XCJC=1 FC=0.170253 CJS=0 VJS=0.75 MJS=0.5 TR=1e-07 PTF=0 KF=0 AF=1)

